`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Module Name: tb_debug_unit
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
// Qu� quiero probar? 
// - Mandar por uart (rx) los comandos para ir pasando de estado,
// ver qu� salidas hay.
// - Poner una memoria (instrucciones) y analizar si puedo pasar el contenido de una memoria a otra por uart
// - Poner banco de registros y ver si esos datos se env�an bien
// - Armar todo lo anterior y probarlo en otro tb con sintesis e implementacion
//////////////////////////////////////////////////////////////////////////////////


module tb_debug_unit(

    );
endmodule
